module malvar_he_cutler_demosaic_tb ();
    malvar_he_cutler_demosaic malvar_he_cutler_demosaic();
    initial
    begin
        $finish;
    end
endmodule
